module ProgramRegister(HBOut, VBOut,AIPOut, AILOut);
output reg[1:0] HBOut=0;
output reg[1:0] VBOut=2;
output reg[3:0] AIPOut=10;
output reg[3:0] AILOut=10;
endmodule
